LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY control_l IS
    PORT (ir     		: IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
			 mode			: IN  STD_LOGIC;
          op     		: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
          ldpc   		: OUT STD_LOGIC;
          wrd    		: OUT STD_LOGIC;
          addr_a 		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			 addr_b 		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
          addr_d 		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
          immed  		: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			 wr_m	  		: OUT STD_LOGIC := '0';
			 in_d			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			 immed_x2	: OUT STD_LOGIC;
			 word_byte	: OUT STD_LOGIC;
			 y_b			: OUT STD_LOGIC;
			 op_salt		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
			 addr_io		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			 wr_out		: OUT STD_LOGIC := '0';
			 rd_in		: OUT STD_LOGIC;
			 a_sys_rd 	: OUT STD_LOGIC;
			 a_sys_wr 	: OUT STD_LOGIC;
			 mask	 	 	: OUT STD_LOGIC;
			 inta			: OUT STD_LOGIC := '0';
			 ilegal_ins : OUT STD_LOGIC := '0';
			 load_store : OUT STD_LOGIC := '0';
			 calls		: OUT STD_LOGIC := '0';
			 mode_exc	: OUT STD_LOGIC := '0';
			 mem_instr	: OUT STD_LOGIC;
			 reti 		: OUT STD_LOGIC := '0');	
END control_l;


ARCHITECTURE Structure OF control_l IS

CONSTANT LOGIC_ARITH	:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT COMPARE		:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
CONSTANT ADDI			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
CONSTANT LOAD			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
CONSTANT STORE			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
CONSTANT MOV			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
CONSTANT BRANCH		:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
CONSTANT IO				:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
CONSTANT MULDIV		: 	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
CONSTANT FLOAT			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
CONSTANT JMP			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
CONSTANT LOADB			:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";
CONSTANT STOREB		:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110";
CONSTANT SYSTEM		:	STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111";


CONSTANT OP_MOVI 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
CONSTANT OP_MOVHI 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
CONSTANT OP_AND 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
CONSTANT OP_OR 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
CONSTANT OP_XOR 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
CONSTANT OP_NOT 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
CONSTANT OP_ADD 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
CONSTANT OP_SUB 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
CONSTANT OP_SHA 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
CONSTANT OP_SHL 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
CONSTANT OP_MUL 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
CONSTANT OP_MULH 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
CONSTANT OP_MULHU 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
CONSTANT OP_DIV 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
CONSTANT OP_DIVU 		:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
CONSTANT OP_CMPLT 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
CONSTANT OP_CMPLE 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
CONSTANT OP_CMPEQ 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
CONSTANT OP_CMPLTU 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
CONSTANT OP_CMPLEU 	:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";

CONSTANT OP_Y			:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "11110"; ----dejamos pasar la y
CONSTANT OP_X			:	STD_LOGIC_VECTOR(4 DOWNTO 0) := "11111"; ----dejamos pasar la x


CONSTANT F_AND			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
CONSTANT F_OR			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
CONSTANT F_XOR			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";
CONSTANT F_NOT			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
CONSTANT F_ADD			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
CONSTANT F_SUB			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";
CONSTANT F_SHA			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
CONSTANT F_SHL			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";

CONSTANT F_CMPLT		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
CONSTANT F_CMPLE		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
CONSTANT F_CMPEQ		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
CONSTANT F_CMPLTU		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
CONSTANT F_CMPLEU		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";

CONSTANT F_MUL			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
CONSTANT F_MULH		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
CONSTANT F_MULHU		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";
CONSTANT F_DIV			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
CONSTANT F_DIVU		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";

CONSTANT F_JZ			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
CONSTANT F_JNZ			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
CONSTANT F_JMP			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
CONSTANT F_JAL			:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
CONSTANT F_CALLS		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";

CONSTANT SYS_RDS		:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "101100";
CONSTANT SYS_WRS		:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "110000";
CONSTANT SYS_EI		:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "100000";
CONSTANT SYS_DI		:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "100001";
CONSTANT SYS_RETI		:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "100100";
CONSTANT SYS_GETIID	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "101000";

CONSTANT SALT_JALJMP	:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";
CONSTANT SALT_JZ		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
CONSTANT SALT_JNZ		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";
CONSTANT SALT_BZ		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
CONSTANT SALT_BNZ		:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
CONSTANT SALT_RETI	:	STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";


SIGNAL HALT		:	STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '1');
SIGNAL EXT		:	STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL OPCODE	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL FCODE	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL SYSCODE	:	STD_LOGIC_VECTOR(5 DOWNTO 0);

--Auxiliars
SIGNAL ldpc_aux			:	STD_LOGIC;
SIGNAL ilegal_ins_aux	: 	STD_LOGIC := '0';

BEGIN
	
	--Auxiliars
	OPCODE <= ir(15 DOWNTO 12);
	
	FCODE  <= 	ir(2 DOWNTO 0) WHEN OPCODE = JMP ELSE
					ir(5 DOWNTO 3);
	
	EXT <= 	(OTHERS => ir(7)) WHEN (OPCODE = MOV OR OPCODE = BRANCH) ELSE	--Extensio de signe segons la operacio
				(OTHERS => ir(5));
				
	SYSCODE	<= ir(5 DOWNTO 0);
	
	--Assignacions output
	
	op <= 	OP_MOVI 		WHEN (OPCODE = MOV 			AND ir(8) = '0') 			ELSE
				OP_MOVHI 	WHEN (OPCODE = MOV 			AND ir(8) = '1') 			ELSE
				OP_AND		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_AND) 		ELSE
				OP_OR			WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_OR) 		ELSE
				OP_XOR		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_XOR) 		ELSE
				OP_NOT		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_NOT) 		ELSE
				OP_ADD		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_ADD) 		ELSE
				OP_SUB		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_SUB) 		ELSE
				OP_SHA		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_SHA) 		ELSE
				OP_SHL		WHEN (OPCODE = LOGIC_ARITH AND FCODE = F_SHL) 		ELSE
				OP_CMPLT		WHEN (OPCODE = COMPARE 		AND FCODE = F_CMPLT) 	ELSE
				OP_CMPLE		WHEN (OPCODE = COMPARE 		AND FCODE = F_CMPLE) 	ELSE
				OP_CMPEQ		WHEN (OPCODE = COMPARE 		AND FCODE = F_CMPEQ) 	ELSE
				OP_CMPLTU	WHEN (OPCODE = COMPARE 		AND FCODE = F_CMPLTU)	ELSE
				OP_CMPLEU	WHEN (OPCODE = COMPARE 		AND FCODE = F_CMPLEU) 	ELSE
				OP_MUL 		WHEN (OPCODE = MULDIV 		AND FCODE = F_MUL) 		ELSE
				OP_MULH 		WHEN (OPCODE = MULDIV 		AND FCODE = F_MULH)		ELSE
				OP_MULHU		WHEN (OPCODE = MULDIV 		AND FCODE = F_MULHU) 	ELSE
				OP_DIV 		WHEN (OPCODE = MULDIV 		AND FCODE = F_DIV) 		ELSE
				OP_DIVU 		WHEN (OPCODE = MULDIV 		AND FCODE = F_DIVU) 		ELSE
				OP_X 			WHEN (OPCODE = SYSTEM 		AND (SYSCODE = SYS_RETI OR 
																	SYSCODE = SYS_RDS  		OR 
																	SYSCODE = SYS_WRS))		ELSE
				OP_Y 			WHEN (OPCODE = SYSTEM 		AND (SYSCODE = SYS_EI 	OR
																	SYSCODE = SYS_DI))		ELSE
				OP_ADD; --inclou ADDI i accessos a memoria
	
	y_b <= 	'0' WHEN (	OPCODE = MOV OR OPCODE = ADDI OR OPCODE = LOAD OR
								OPCODE = STORE OR OPCODE = LOADB OR OPCODE = STOREB
								OR (OPCODE = SYSTEM AND (SYSCODE = SYS_EI OR
																	SYSCODE = SYS_DI))) ELSE
				'1';
	
	ldpc_aux <= 	'0' WHEN ir = HALT ELSE 
						'1';
				
	ldpc <= ldpc_aux;			
	
	wrd <= 	'0' WHEN (ilegal_ins_aux = '1') ELSE	-- If ilegal instruction, no write permission
				'1' WHEN (ldpc_aux = '1' AND (	OPCODE = LOGIC_ARITH OR 
															OPCODE = LOAD			OR
															OPCODE = MOV			OR
															OPCODE = LOADB			OR
															OPCODE = ADDI			OR
															OPCODE = MULDIV		OR
															OPCODE = COMPARE		OR
															OPCODE = SYSTEM		OR
															(OPCODE = JMP AND (FCODE = F_JAL OR FCODE = F_CALLS)) OR
															(OPCODE = IO AND ir(8) = '0'))) 	ELSE
				'0';
	
	addr_a <= 	"000"					WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_RETI)	ELSE
					ir(11 DOWNTO 9) 	WHEN (OPCODE = MOV)										ELSE
					ir(8 DOWNTO 6);
	
	addr_b <= 	"001"					WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_RETI)	ELSE
					ir(2 DOWNTO 0) 	WHEN (OPCODE = LOGIC_ARITH OR OPCODE = COMPARE OR OPCODE = MULDIV) 	ELSE
					ir(11 DOWNTO 9);
					
	addr_d <= 	"111"					WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_RETI)	ELSE
					"011"					WHEN (OPCODE = JMP 	 AND FCODE = F_CALLS)		ELSE
					ir(11 DOWNTO 9);
	
	immed <= "0000000000000001"	WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_EI)			ELSE
				"0000000000000000"	WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_DI)			ELSE
				EXT(7 DOWNTO 0) & ir(7 DOWNTO 0) WHEN (OPCODE = MOV OR OPCODE = BRANCH) ELSE
				EXT & ir(5 DOWNTO 0);
	
	wr_m <= 	'1' WHEN (OPCODE = STORE OR OPCODE = STOREB) AND (ilegal_ins_aux = '0') ELSE	--Store, Load AND no ilegal ins.
				'0';
	
	in_d <= 	"011" WHEN ((OPCODE = IO AND ir(8) = '0') OR
							  (OPCODE = SYSTEM AND SYSCODE = SYS_GETIID)) 	ELSE
				"010" WHEN (OPCODE = JMP AND FCODE = F_JAL) 					ELSE
				"001" WHEN (OPCODE = LOAD OR OPCODE = LOADB) 				ELSE
				"000";
	 
	immed_x2 <= 	'1' WHEN (OPCODE = LOAD OR OPCODE = STORE OR OPCODE = BRANCH) ELSE
						'0';
	
	word_byte <= 	'1' WHEN (OPCODE = LOADB OR OPCODE = STOREB) ELSE
						'0';
						
	op_salt <=	"000"			WHEN ilegal_ins_aux = '1'													ELSE 	-- When the instruction doesn't exist, no jump.
					SALT_JALJMP	WHEN (OPCODE = JMP AND (FCODE = F_JAL OR FCODE = F_JMP))			ELSE --Inconditional jumps
					SALT_JZ		WHEN (OPCODE = JMP AND (FCODE = F_JZ))									ELSE --Rest of jumps JZ
					SALT_JNZ 	WHEN (OPCODE = JMP AND (FCODE = F_JNZ))								ELSE --Rest of jumps JNZ
					SALT_BZ		WHEN (OPCODE = BRANCH AND ir(8) = '0')									ELSE --Branchs BZ
					SALT_BNZ 	WHEN (OPCODE = BRANCH AND ir(8) = '1')									ELSE --Branchs BNZ
					SALT_RETI	WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_RETI AND mode = '1')	ELSE --RETI
					"000";	--Rest of operations
				
	addr_io	<= ir(7 DOWNTO 0);
	
	wr_out <= 	'1' WHEN OPCODE = IO AND ir(8) = '1' AND ilegal_ins_aux = '0' ELSE
					'0';
				
	rd_in  <= 	'1' WHEN ((OPCODE = IO AND ir(8) = '0') OR
								(OPCODE = SYSTEM AND SYSCODE = SYS_GETIID)) ELSE
					'0';
	
	a_sys_rd	<= '1' WHEN (OPCODE = SYSTEM AND (	SYSCODE = SYS_RETI 	OR
																SYSCODE = SYS_RDS))		ELSE
					'0';
					
	a_sys_wr	<= '1' WHEN (	(OPCODE = JMP 	 AND FCODE = F_CALLS)		OR
									(OPCODE = SYSTEM AND (SYSCODE = SYS_WRS 	OR
																SYSCODE = SYS_EI		OR
																SYSCODE = SYS_DI		OR
																SYSCODE = SYS_RETI)))		ELSE
					'0';
					
	mask	<= '1' WHEN (OPCODE = SYSTEM AND (	SYSCODE = SYS_EI 	OR
															SYSCODE = SYS_DI))			ELSE
				'0';
				
	inta <= 	'1' 	WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_GETIID AND ilegal_ins_aux = '0') ELSE
				'0';		
				
	ilegal_ins_aux <=  '1' WHEN (	(OPCODE = COMPARE AND FCODE = "010") 				OR
										(OPCODE = COMPARE AND FCODE = "110") 					OR
										(OPCODE = COMPARE AND FCODE = "111") 					OR
										(OPCODE = MULDIV  AND FCODE = "011") 					OR
										(OPCODE = MULDIV  AND FCODE = "110") 					OR
										(OPCODE = MULDIV  AND FCODE = "111") 					OR	
										(OPCODE = FLOAT)												OR
										(OPCODE = JMP AND ir(5 DOWNTO 3) /= "000") 			OR
										(OPCODE = JMP AND (FCODE = F_JMP OR FCODE = F_CALLS) AND ir(11 DOWNTO 9) /= "000") OR
										(OPCODE = JMP AND FCODE = F_CALLS AND mode = '1') 	OR	--Calls en modo sistema
										(OPCODE = JMP AND FCODE = "010") 						OR
										(OPCODE = JMP AND FCODE = "101") 						OR
										(OPCODE = JMP AND FCODE = "110") 						OR
										(OPCODE = SYSTEM AND ir(5) = '0') 						OR
										(OPCODE = SYSTEM AND (	SYSCODE /= SYS_RDS 			AND
																		SYSCODE /= SYS_WRS 			AND
																		SYSCODE /= SYS_EI	 			AND
																		SYSCODE /= SYS_DI	 			AND
																		SYSCODE /= SYS_RETI 			AND
																		SYSCODE /= SYS_GETIID		AND
																		ir /= HALT)) 					OR
										(OPCODE = SYSTEM AND (SYSCODE = SYS_EI OR SYSCODE = SYS_DI OR SYSCODE = SYS_RETI) AND ir(11 DOWNTO 6) /= "000000") OR
										(OPCODE = SYSTEM AND SYSCODE = SYS_GETIID AND ir(8 DOWNTO 6) /= "000")) ELSE			
						'0';
						
	ilegal_ins <= ilegal_ins_aux;

	load_store <= 	'1' WHEN 	(OPCODE = LOAD OR OPCODE = STORE)	ELSE
						'0';

	calls <=	'1' WHEN (OPCODE = JMP AND FCODE = F_CALLS)	ELSE
				'0';
				
	--Trying to execute a system instruction while on user mode.
	mode_exc	<=	'1' WHEN (OPCODE = SYSTEM AND mode = '0' AND (	SYSCODE = SYS_RDS 	OR
																					SYSCODE = SYS_WRS 	OR
																					SYSCODE = SYS_EI	 	OR
																					SYSCODE = SYS_DI	 	OR
																					SYSCODE = SYS_RETI 	OR
																					SYSCODE = SYS_GETIID )	) ELSE
					'0';
					
	mem_instr <= 	'1' WHEN (OPCODE = LOAD OR OPCODE = STORE OR OPCODE = LOADB OR OPCODE = STOREB) ELSE
						'0';
	
	reti <=	'1' WHEN (OPCODE = SYSTEM AND SYSCODE = SYS_RETI) ELSE
				'0';
	
END Structure;